/******************************
made 2019/1/30 powered harumaki
module name: activation
this is activation function

only ReLU
*******************************/

module activation();
    
endmodule