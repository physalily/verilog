/******************************
made 2019/1/25 powered harumaki
module name: CoreSocket
this is 

function list
*******************************/

module CoreSocket();

    begin
    MatrixCore(
        
        );
    end
endmodule