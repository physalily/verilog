/******************************
made 2019/2/3 powered harumaki
module name: inst_decoder
this is instruction decoder
function list
*******************************/

module inst_decoder();
    
endmodule